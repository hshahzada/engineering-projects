library verilog;
use verilog.vl_types.all;
entity decodmodified_vlg_vec_tst is
end decodmodified_vlg_vec_tst;
