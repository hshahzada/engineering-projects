library verilog;
use verilog.vl_types.all;
entity johns_vlg_vec_tst is
end johns_vlg_vec_tst;
