library verilog;
use verilog.vl_types.all;
entity C_vlg_vec_tst is
end C_vlg_vec_tst;
